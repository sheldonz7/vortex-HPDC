// this is a temporary file we can use for the vortex adapter