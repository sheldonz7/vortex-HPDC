// this is a temporary file we can use for the vortex adapter

// in the cva6 repo, this file served the purpose of mapping its core’s request and response signals to the HPDCache

//THINGS WE NEED:
// * handle input output requests
// * Atomic operations? (these were included in cva6 and I am not quite sure if they are needed here)
// * Flush mannagement? (these were included in cva6 and I am not quite sure if they are needed here)
// * possible bank routing and mannagement 